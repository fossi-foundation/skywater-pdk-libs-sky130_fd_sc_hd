# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.370000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.085000  0.085000 0.375000 0.810000 ;
        RECT 2.020000  0.085000 2.350000 0.895000 ;
        RECT 3.115000  0.085000 3.445000 0.900000 ;
        RECT 3.975000  0.085000 4.305000 0.560000 ;
        RECT 4.835000  0.085000 5.165000 0.900000 ;
        RECT 5.825000  0.085000 6.155000 0.900000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000000 5.355000 6.440000 5.525000 ;
        RECT 0.085000 4.630000 0.375000 5.355000 ;
        RECT 2.645000 4.515000 2.905000 5.355000 ;
        RECT 3.575000 4.515000 3.765000 5.355000 ;
        RECT 4.445000 4.515000 4.955000 5.355000 ;
        RECT 6.065000 4.630000 6.355000 5.355000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.890000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.890000 1.625000 5.120000 2.635000 ;
        RECT 4.890000 2.635000 6.440000 2.805000 ;
        RECT 4.890000 2.805000 5.120000 3.740000 ;
        RECT 5.905000 1.610000 6.075000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.560000 0.375000 2.800000 2.130000 ;
      RECT 2.560000 2.130000 3.390000 2.370000 ;
      RECT 3.060000 2.370000 3.390000 3.965000 ;
      RECT 3.075000 4.265000 4.265000 4.325000 ;
      RECT 3.075000 4.325000 3.405000 5.185000 ;
      RECT 3.145000 4.155000 4.195000 4.265000 ;
      RECT 3.615000 0.255000 3.805000 0.730000 ;
      RECT 3.615000 0.730000 4.665000 0.980000 ;
      RECT 3.680000 2.405000 4.190000 2.575000 ;
      RECT 3.680000 2.575000 3.850000 3.470000 ;
      RECT 3.680000 3.470000 4.720000 3.640000 ;
      RECT 3.935000 4.325000 4.265000 5.185000 ;
      RECT 4.020000 0.980000 4.190000 2.405000 ;
      RECT 4.020000 2.745000 4.640000 2.915000 ;
      RECT 4.020000 2.915000 4.190000 3.300000 ;
      RECT 4.020000 3.810000 4.190000 4.155000 ;
      RECT 4.390000 3.085000 4.720000 3.470000 ;
      RECT 4.410000 3.640000 4.720000 3.740000 ;
      RECT 4.470000 1.625000 4.640000 2.745000 ;
      RECT 4.475000 0.255000 4.665000 0.730000 ;
      RECT 5.135000 4.405000 5.765000 4.460000 ;
      RECT 5.135000 4.460000 5.695000 4.820000 ;
      RECT 5.135000 4.820000 5.485000 5.160000 ;
      RECT 5.360000 3.070000 5.550000 4.125000 ;
      RECT 5.360000 4.125000 6.085000 4.355000 ;
      RECT 5.360000 4.355000 5.765000 4.405000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
END LIBRARY
